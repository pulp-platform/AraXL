// Copyright 2021-2025 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Author: Matheus Cavalcante <matheusd@iis.ee.ethz.ch>
// Date: 21/10/2020
// Description: Top level testbench module for Verilator.

module ara_tb_verilator #(
    parameter int unsigned NrLanes = 0,
    parameter int unsigned NrClusters = 0
  )(
    input  logic        clk_i,
    input  logic        rst_ni,
    output logic [63:0] exit_o
  );

  /*****************
   *  Definitions  *
   *****************/

  // localparam AxiAddrWidth     = 64;
  // localparam AxiWideDataWidth = 64 * NrLanes / 2;
  localparam AxiAddrWidth          = 64;
  localparam AxiWideDataWidth      = 32 * NrLanes * NrClusters;
  localparam ClusterAxiDataWidth   = 32 * NrLanes;

  /*********
   *  DUT  *
   *********/

  // ara_testharness #(
  //   .NrLanes     (NrLanes         ),
  //   .AxiAddrWidth(AxiAddrWidth    ),
  //   .AxiDataWidth(AxiWideDataWidth)
  // ) dut (
  //   .clk_i (clk_i ),
  //   .rst_ni(rst_ni),
  //   .exit_o(exit_o)
  // );

  ara_testharness #(
    .NrLanes     (NrLanes         ),
    .NrClusters  (NrClusters      ),
    .AxiAddrWidth(AxiAddrWidth    ),
    .AxiDataWidth(AxiWideDataWidth),
    .ClusterAxiDataWidth(ClusterAxiDataWidth)
  ) dut (
    .clk_i (clk_i ),
    .rst_ni(rst_ni),
    .exit_o(exit_o)
  );

  /*********
   *  EOC  *
   *********/

  always @(posedge clk_i) begin
    if (exit_o[0]) begin
      if (exit_o >> 1) begin
        $warning("Core Test ", $sformatf("*** FAILED *** (tohost = %0d)", (exit_o >> 1)));
      end else begin
        // Print vector HW runtime
        $display("[hw-cycles]: %d", int'(dut.runtime_buf_q));
        $info("Core Test ", $sformatf("*** SUCCESS *** (tohost = %0d)", (exit_o >> 1)));
      end

      $finish(exit_o >> 1);
    end
  end

endmodule : ara_tb_verilator
