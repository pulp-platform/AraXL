// Copyright 2023-2025 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Author: Matteo Perotti <mperotti@iis.ee.ethz.ch>
// Description:
// Ara's optimized SLDU datapath.
// Cannot reshuffle AND slide at the same time.

module sldu_op_dp import ara_pkg::*; import rvv_pkg::*; import cf_math_pkg::idx_width; #(
    parameter int unsigned NrLanes = 0,
    // Dependant parameters. DO NOT CHANGE!
    localparam int  unsigned DataWidth = $bits(elen_t), // Width of the lane datapath
    localparam int  unsigned StrbWidth = DataWidth/8,
    localparam type          strb_t    = logic [StrbWidth-1:0] // Byte-strobe type
  ) (
    input  elen_t                      [NrLanes-1:0] op_i,
    input  logic            [idx_width(4*NrLanes):0] slamt_i,
    input  rvv_pkg::vew_e                            eew_src_i,
    input  rvv_pkg::vew_e                            eew_dst_i,
    input  logic                                     dir_i,
    output elen_t                      [NrLanes-1:0] op_o
);

logic [$bits(op_i)-1:0] op_i_flat;
logic [$bits(op_o)-1:0] op_o_flat;

assign op_i_flat = op_i;
assign op_o      = op_o_flat;

if (NrLanes == 1)
  always_comb begin
    unique case ({eew_src_i, eew_dst_i, slamt_i, dir_i})
      {EW8, EW8, 3'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW8, EW16, 3'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW8, EW32, 3'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW8, EW64, 3'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW8, EW8, 3'd1, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[24 +: 8];
      end
      {EW8, EW8, 3'd1, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[0 +: 8];
      end
      {EW8, EW8, 3'd2, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[40 +: 8];
      end
      {EW8, EW8, 3'd2, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[32 +: 8];
      end
      {EW8, EW8, 3'd4, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[48 +: 8];
      end
      {EW8, EW8, 3'd4, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[48 +: 8];
      end
      {EW16, EW8, 3'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW16, EW16, 3'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW16, EW32, 3'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW16, EW64, 3'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW16, EW16, 3'd1, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[24 +: 8];
      end
      {EW16, EW16, 3'd1, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[8 +: 8];
      end
      {EW16, EW16, 3'd2, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[40 +: 8];
      end
      {EW16, EW16, 3'd2, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[40 +: 8];
      end
      {EW16, EW16, 3'd4, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW16, EW16, 3'd4, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW32, EW8, 3'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW32, EW16, 3'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW32, EW32, 3'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW32, EW64, 3'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW32, EW32, 3'd1, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[24 +: 8];
      end
      {EW32, EW32, 3'd1, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[24 +: 8];
      end
      {EW32, EW32, 3'd2, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW32, EW32, 3'd2, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW32, EW32, 3'd4, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW32, EW32, 3'd4, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW64, EW8, 3'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW64, EW16, 3'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW64, EW32, 3'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW64, EW64, 3'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW64, EW64, 3'd1, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW64, EW64, 3'd1, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW64, EW64, 3'd2, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW64, EW64, 3'd2, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW64, EW64, 3'd4, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      {EW64, EW64, 3'd4, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
      end
      default: op_o_flat = op_i_flat;
    endcase
  end
else if (NrLanes == 2)
  always_comb begin
    unique case ({eew_src_i, eew_dst_i, slamt_i, dir_i})
      {EW8, EW8, 4'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW8, EW16, 4'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW8, EW32, 4'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW8, EW64, 4'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW8, EW8, 4'd1, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[56 +: 8];
      end
      {EW8, EW8, 4'd1, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[0 +: 8];
      end
      {EW8, EW8, 4'd2, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[88 +: 8];
      end
      {EW8, EW8, 4'd2, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[64 +: 8];
      end
      {EW8, EW8, 4'd4, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[104 +: 8];
      end
      {EW8, EW8, 4'd4, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[96 +: 8];
      end
      {EW8, EW8, 4'd8, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[112 +: 8];
      end
      {EW8, EW8, 4'd8, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[112 +: 8];
      end
      {EW16, EW8, 4'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW16, EW16, 4'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW16, EW32, 4'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW16, EW64, 4'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW16, EW16, 4'd1, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[56 +: 8];
      end
      {EW16, EW16, 4'd1, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[8 +: 8];
      end
      {EW16, EW16, 4'd2, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[88 +: 8];
      end
      {EW16, EW16, 4'd2, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[72 +: 8];
      end
      {EW16, EW16, 4'd4, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[104 +: 8];
      end
      {EW16, EW16, 4'd4, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[104 +: 8];
      end
      {EW16, EW16, 4'd8, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW16, EW16, 4'd8, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW32, EW8, 4'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW32, EW16, 4'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW32, EW32, 4'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW32, EW64, 4'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW32, EW32, 4'd1, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[56 +: 8];
      end
      {EW32, EW32, 4'd1, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[24 +: 8];
      end
      {EW32, EW32, 4'd2, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[88 +: 8];
      end
      {EW32, EW32, 4'd2, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[88 +: 8];
      end
      {EW32, EW32, 4'd4, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW32, EW32, 4'd4, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW32, EW32, 4'd8, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW32, EW32, 4'd8, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW64, EW8, 4'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW64, EW16, 4'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW64, EW32, 4'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW64, EW64, 4'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW64, EW64, 4'd1, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[56 +: 8];
      end
      {EW64, EW64, 4'd1, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[56 +: 8];
      end
      {EW64, EW64, 4'd2, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW64, EW64, 4'd2, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW64, EW64, 4'd4, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW64, EW64, 4'd4, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW64, EW64, 4'd8, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      {EW64, EW64, 4'd8, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
      end
      default: op_o_flat = op_i_flat;
    endcase
  end
else if (NrLanes == 4)
  always_comb begin
    unique case ({eew_src_i, eew_dst_i, slamt_i, dir_i})
      {EW8, EW8, 5'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW8, EW16, 5'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW8, EW32, 5'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW8, EW64, 5'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW8, EW8, 5'd1, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[184 +: 8];
      end
      {EW8, EW8, 5'd1, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[0 +: 8];
      end
      {EW8, EW8, 5'd2, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[120 +: 8];
      end
      {EW8, EW8, 5'd2, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[64 +: 8];
      end
      {EW8, EW8, 5'd4, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[216 +: 8];
      end
      {EW8, EW8, 5'd4, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[192 +: 8];
      end
      {EW8, EW8, 5'd8, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[232 +: 8];
      end
      {EW8, EW8, 5'd8, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[224 +: 8];
      end
      {EW8, EW8, 5'd16, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[240 +: 8];
      end
      {EW8, EW8, 5'd16, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[240 +: 8];
      end
      {EW16, EW8, 5'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW16, EW16, 5'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW16, EW32, 5'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW16, EW64, 5'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW16, EW16, 5'd1, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[184 +: 8];
      end
      {EW16, EW16, 5'd1, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[8 +: 8];
      end
      {EW16, EW16, 5'd2, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[120 +: 8];
      end
      {EW16, EW16, 5'd2, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[72 +: 8];
      end
      {EW16, EW16, 5'd4, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[216 +: 8];
      end
      {EW16, EW16, 5'd4, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[200 +: 8];
      end
      {EW16, EW16, 5'd8, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[232 +: 8];
      end
      {EW16, EW16, 5'd8, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[232 +: 8];
      end
      {EW16, EW16, 5'd16, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW16, EW16, 5'd16, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW32, EW8, 5'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW32, EW16, 5'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW32, EW32, 5'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW32, EW64, 5'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW32, EW32, 5'd1, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[184 +: 8];
      end
      {EW32, EW32, 5'd1, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[24 +: 8];
      end
      {EW32, EW32, 5'd2, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[120 +: 8];
      end
      {EW32, EW32, 5'd2, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[88 +: 8];
      end
      {EW32, EW32, 5'd4, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[216 +: 8];
      end
      {EW32, EW32, 5'd4, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[216 +: 8];
      end
      {EW32, EW32, 5'd8, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW32, EW32, 5'd8, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW32, EW32, 5'd16, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW32, EW32, 5'd16, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW64, EW8, 5'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW64, EW16, 5'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW64, EW32, 5'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW64, EW64, 5'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW64, EW64, 5'd1, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[184 +: 8];
      end
      {EW64, EW64, 5'd1, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[56 +: 8];
      end
      {EW64, EW64, 5'd2, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[120 +: 8];
      end
      {EW64, EW64, 5'd2, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[120 +: 8];
      end
      {EW64, EW64, 5'd4, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW64, EW64, 5'd4, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW64, EW64, 5'd8, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW64, EW64, 5'd8, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW64, EW64, 5'd16, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      {EW64, EW64, 5'd16, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
      end
      default: op_o_flat = op_i_flat;
    endcase
  end
else if (NrLanes == 8)
  always_comb begin
    unique case ({eew_src_i, eew_dst_i, slamt_i, dir_i})
      {EW8, EW8, 6'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW8, EW16, 6'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW8, EW32, 6'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW8, EW64, 6'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW8, EW8, 6'd1, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[440 +: 8];
      end
      {EW8, EW8, 6'd1, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[0 +: 8];
      end
      {EW8, EW8, 6'd2, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[376 +: 8];
      end
      {EW8, EW8, 6'd2, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[64 +: 8];
      end
      {EW8, EW8, 6'd4, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[248 +: 8];
      end
      {EW8, EW8, 6'd4, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[192 +: 8];
      end
      {EW8, EW8, 6'd8, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[472 +: 8];
      end
      {EW8, EW8, 6'd8, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[448 +: 8];
      end
      {EW8, EW8, 6'd16, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[488 +: 8];
      end
      {EW8, EW8, 6'd16, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[480 +: 8];
      end
      {EW8, EW8, 6'd32, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[496 +: 8];
      end
      {EW8, EW8, 6'd32, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[496 +: 8];
      end
      {EW16, EW8, 6'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW16, EW16, 6'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW16, EW32, 6'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW16, EW64, 6'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW16, EW16, 6'd1, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[440 +: 8];
      end
      {EW16, EW16, 6'd1, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[8 +: 8];
      end
      {EW16, EW16, 6'd2, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[376 +: 8];
      end
      {EW16, EW16, 6'd2, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[72 +: 8];
      end
      {EW16, EW16, 6'd4, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[248 +: 8];
      end
      {EW16, EW16, 6'd4, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[200 +: 8];
      end
      {EW16, EW16, 6'd8, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[472 +: 8];
      end
      {EW16, EW16, 6'd8, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[456 +: 8];
      end
      {EW16, EW16, 6'd16, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[488 +: 8];
      end
      {EW16, EW16, 6'd16, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[488 +: 8];
      end
      {EW16, EW16, 6'd32, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW16, EW16, 6'd32, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW32, EW8, 6'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW32, EW16, 6'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW32, EW32, 6'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW32, EW64, 6'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW32, EW32, 6'd1, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[440 +: 8];
      end
      {EW32, EW32, 6'd1, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[24 +: 8];
      end
      {EW32, EW32, 6'd2, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[376 +: 8];
      end
      {EW32, EW32, 6'd2, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[88 +: 8];
      end
      {EW32, EW32, 6'd4, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[248 +: 8];
      end
      {EW32, EW32, 6'd4, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[216 +: 8];
      end
      {EW32, EW32, 6'd8, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[472 +: 8];
      end
      {EW32, EW32, 6'd8, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[472 +: 8];
      end
      {EW32, EW32, 6'd16, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW32, EW32, 6'd16, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW32, EW32, 6'd32, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW32, EW32, 6'd32, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW64, EW8, 6'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW64, EW16, 6'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW64, EW32, 6'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW64, EW64, 6'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW64, EW64, 6'd1, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[440 +: 8];
      end
      {EW64, EW64, 6'd1, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[56 +: 8];
      end
      {EW64, EW64, 6'd2, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[376 +: 8];
      end
      {EW64, EW64, 6'd2, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[120 +: 8];
      end
      {EW64, EW64, 6'd4, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[248 +: 8];
      end
      {EW64, EW64, 6'd4, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[248 +: 8];
      end
      {EW64, EW64, 6'd8, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW64, EW64, 6'd8, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW64, EW64, 6'd16, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW64, EW64, 6'd16, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW64, EW64, 6'd32, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      {EW64, EW64, 6'd32, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
      end
      default: op_o_flat = op_i_flat;
    endcase
  end
else if (NrLanes == 16)
  always_comb begin
    unique case ({eew_src_i, eew_dst_i, slamt_i, dir_i})
      {EW8, EW8, 7'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW8, EW16, 7'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW8, EW32, 7'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW8, EW64, 7'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW8, EW8, 7'd1, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[952 +: 8];
      end
      {EW8, EW8, 7'd1, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[0 +: 8];
      end
      {EW8, EW8, 7'd2, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[888 +: 8];
      end
      {EW8, EW8, 7'd2, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[64 +: 8];
      end
      {EW8, EW8, 7'd4, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[760 +: 8];
      end
      {EW8, EW8, 7'd4, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[192 +: 8];
      end
      {EW8, EW8, 7'd8, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[504 +: 8];
      end
      {EW8, EW8, 7'd8, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[448 +: 8];
      end
      {EW8, EW8, 7'd16, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[984 +: 8];
      end
      {EW8, EW8, 7'd16, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[960 +: 8];
      end
      {EW8, EW8, 7'd32, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1000 +: 8];
      end
      {EW8, EW8, 7'd32, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[992 +: 8];
      end
      {EW8, EW8, 7'd64, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1008 +: 8];
      end
      {EW8, EW8, 7'd64, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1008 +: 8];
      end
      {EW16, EW8, 7'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW16, EW16, 7'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW16, EW32, 7'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW16, EW64, 7'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW16, EW16, 7'd1, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[952 +: 8];
      end
      {EW16, EW16, 7'd1, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[8 +: 8];
      end
      {EW16, EW16, 7'd2, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[888 +: 8];
      end
      {EW16, EW16, 7'd2, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[72 +: 8];
      end
      {EW16, EW16, 7'd4, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[760 +: 8];
      end
      {EW16, EW16, 7'd4, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[200 +: 8];
      end
      {EW16, EW16, 7'd8, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[504 +: 8];
      end
      {EW16, EW16, 7'd8, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[456 +: 8];
      end
      {EW16, EW16, 7'd16, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[984 +: 8];
      end
      {EW16, EW16, 7'd16, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[968 +: 8];
      end
      {EW16, EW16, 7'd32, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1000 +: 8];
      end
      {EW16, EW16, 7'd32, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1000 +: 8];
      end
      {EW16, EW16, 7'd64, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW16, EW16, 7'd64, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW32, EW8, 7'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW32, EW16, 7'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW32, EW32, 7'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW32, EW64, 7'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW32, EW32, 7'd1, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[952 +: 8];
      end
      {EW32, EW32, 7'd1, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[24 +: 8];
      end
      {EW32, EW32, 7'd2, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[888 +: 8];
      end
      {EW32, EW32, 7'd2, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[88 +: 8];
      end
      {EW32, EW32, 7'd4, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[760 +: 8];
      end
      {EW32, EW32, 7'd4, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[216 +: 8];
      end
      {EW32, EW32, 7'd8, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[504 +: 8];
      end
      {EW32, EW32, 7'd8, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[472 +: 8];
      end
      {EW32, EW32, 7'd16, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[984 +: 8];
      end
      {EW32, EW32, 7'd16, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[984 +: 8];
      end
      {EW32, EW32, 7'd32, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW32, EW32, 7'd32, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW32, EW32, 7'd64, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW32, EW32, 7'd64, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW64, EW8, 7'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW64, EW16, 7'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW64, EW32, 7'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW64, EW64, 7'd0, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW64, EW64, 7'd1, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[952 +: 8];
      end
      {EW64, EW64, 7'd1, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[56 +: 8];
      end
      {EW64, EW64, 7'd2, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[888 +: 8];
      end
      {EW64, EW64, 7'd2, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[120 +: 8];
      end
      {EW64, EW64, 7'd4, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[760 +: 8];
      end
      {EW64, EW64, 7'd4, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[248 +: 8];
      end
      {EW64, EW64, 7'd8, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[504 +: 8];
      end
      {EW64, EW64, 7'd8, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[1016 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[504 +: 8];
      end
      {EW64, EW64, 7'd16, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW64, EW64, 7'd16, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW64, EW64, 7'd32, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW64, EW64, 7'd32, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW64, EW64, 7'd64, 1'b1}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      {EW64, EW64, 7'd64, 1'b0}: begin
        op_o_flat[0 +: 8] = op_i_flat[0 +: 8];
        op_o_flat[8 +: 8] = op_i_flat[8 +: 8];
        op_o_flat[16 +: 8] = op_i_flat[16 +: 8];
        op_o_flat[24 +: 8] = op_i_flat[24 +: 8];
        op_o_flat[32 +: 8] = op_i_flat[32 +: 8];
        op_o_flat[40 +: 8] = op_i_flat[40 +: 8];
        op_o_flat[48 +: 8] = op_i_flat[48 +: 8];
        op_o_flat[56 +: 8] = op_i_flat[56 +: 8];
        op_o_flat[64 +: 8] = op_i_flat[64 +: 8];
        op_o_flat[72 +: 8] = op_i_flat[72 +: 8];
        op_o_flat[80 +: 8] = op_i_flat[80 +: 8];
        op_o_flat[88 +: 8] = op_i_flat[88 +: 8];
        op_o_flat[96 +: 8] = op_i_flat[96 +: 8];
        op_o_flat[104 +: 8] = op_i_flat[104 +: 8];
        op_o_flat[112 +: 8] = op_i_flat[112 +: 8];
        op_o_flat[120 +: 8] = op_i_flat[120 +: 8];
        op_o_flat[128 +: 8] = op_i_flat[128 +: 8];
        op_o_flat[136 +: 8] = op_i_flat[136 +: 8];
        op_o_flat[144 +: 8] = op_i_flat[144 +: 8];
        op_o_flat[152 +: 8] = op_i_flat[152 +: 8];
        op_o_flat[160 +: 8] = op_i_flat[160 +: 8];
        op_o_flat[168 +: 8] = op_i_flat[168 +: 8];
        op_o_flat[176 +: 8] = op_i_flat[176 +: 8];
        op_o_flat[184 +: 8] = op_i_flat[184 +: 8];
        op_o_flat[192 +: 8] = op_i_flat[192 +: 8];
        op_o_flat[200 +: 8] = op_i_flat[200 +: 8];
        op_o_flat[208 +: 8] = op_i_flat[208 +: 8];
        op_o_flat[216 +: 8] = op_i_flat[216 +: 8];
        op_o_flat[224 +: 8] = op_i_flat[224 +: 8];
        op_o_flat[232 +: 8] = op_i_flat[232 +: 8];
        op_o_flat[240 +: 8] = op_i_flat[240 +: 8];
        op_o_flat[248 +: 8] = op_i_flat[248 +: 8];
        op_o_flat[256 +: 8] = op_i_flat[256 +: 8];
        op_o_flat[264 +: 8] = op_i_flat[264 +: 8];
        op_o_flat[272 +: 8] = op_i_flat[272 +: 8];
        op_o_flat[280 +: 8] = op_i_flat[280 +: 8];
        op_o_flat[288 +: 8] = op_i_flat[288 +: 8];
        op_o_flat[296 +: 8] = op_i_flat[296 +: 8];
        op_o_flat[304 +: 8] = op_i_flat[304 +: 8];
        op_o_flat[312 +: 8] = op_i_flat[312 +: 8];
        op_o_flat[320 +: 8] = op_i_flat[320 +: 8];
        op_o_flat[328 +: 8] = op_i_flat[328 +: 8];
        op_o_flat[336 +: 8] = op_i_flat[336 +: 8];
        op_o_flat[344 +: 8] = op_i_flat[344 +: 8];
        op_o_flat[352 +: 8] = op_i_flat[352 +: 8];
        op_o_flat[360 +: 8] = op_i_flat[360 +: 8];
        op_o_flat[368 +: 8] = op_i_flat[368 +: 8];
        op_o_flat[376 +: 8] = op_i_flat[376 +: 8];
        op_o_flat[384 +: 8] = op_i_flat[384 +: 8];
        op_o_flat[392 +: 8] = op_i_flat[392 +: 8];
        op_o_flat[400 +: 8] = op_i_flat[400 +: 8];
        op_o_flat[408 +: 8] = op_i_flat[408 +: 8];
        op_o_flat[416 +: 8] = op_i_flat[416 +: 8];
        op_o_flat[424 +: 8] = op_i_flat[424 +: 8];
        op_o_flat[432 +: 8] = op_i_flat[432 +: 8];
        op_o_flat[440 +: 8] = op_i_flat[440 +: 8];
        op_o_flat[448 +: 8] = op_i_flat[448 +: 8];
        op_o_flat[456 +: 8] = op_i_flat[456 +: 8];
        op_o_flat[464 +: 8] = op_i_flat[464 +: 8];
        op_o_flat[472 +: 8] = op_i_flat[472 +: 8];
        op_o_flat[480 +: 8] = op_i_flat[480 +: 8];
        op_o_flat[488 +: 8] = op_i_flat[488 +: 8];
        op_o_flat[496 +: 8] = op_i_flat[496 +: 8];
        op_o_flat[504 +: 8] = op_i_flat[504 +: 8];
        op_o_flat[512 +: 8] = op_i_flat[512 +: 8];
        op_o_flat[520 +: 8] = op_i_flat[520 +: 8];
        op_o_flat[528 +: 8] = op_i_flat[528 +: 8];
        op_o_flat[536 +: 8] = op_i_flat[536 +: 8];
        op_o_flat[544 +: 8] = op_i_flat[544 +: 8];
        op_o_flat[552 +: 8] = op_i_flat[552 +: 8];
        op_o_flat[560 +: 8] = op_i_flat[560 +: 8];
        op_o_flat[568 +: 8] = op_i_flat[568 +: 8];
        op_o_flat[576 +: 8] = op_i_flat[576 +: 8];
        op_o_flat[584 +: 8] = op_i_flat[584 +: 8];
        op_o_flat[592 +: 8] = op_i_flat[592 +: 8];
        op_o_flat[600 +: 8] = op_i_flat[600 +: 8];
        op_o_flat[608 +: 8] = op_i_flat[608 +: 8];
        op_o_flat[616 +: 8] = op_i_flat[616 +: 8];
        op_o_flat[624 +: 8] = op_i_flat[624 +: 8];
        op_o_flat[632 +: 8] = op_i_flat[632 +: 8];
        op_o_flat[640 +: 8] = op_i_flat[640 +: 8];
        op_o_flat[648 +: 8] = op_i_flat[648 +: 8];
        op_o_flat[656 +: 8] = op_i_flat[656 +: 8];
        op_o_flat[664 +: 8] = op_i_flat[664 +: 8];
        op_o_flat[672 +: 8] = op_i_flat[672 +: 8];
        op_o_flat[680 +: 8] = op_i_flat[680 +: 8];
        op_o_flat[688 +: 8] = op_i_flat[688 +: 8];
        op_o_flat[696 +: 8] = op_i_flat[696 +: 8];
        op_o_flat[704 +: 8] = op_i_flat[704 +: 8];
        op_o_flat[712 +: 8] = op_i_flat[712 +: 8];
        op_o_flat[720 +: 8] = op_i_flat[720 +: 8];
        op_o_flat[728 +: 8] = op_i_flat[728 +: 8];
        op_o_flat[736 +: 8] = op_i_flat[736 +: 8];
        op_o_flat[744 +: 8] = op_i_flat[744 +: 8];
        op_o_flat[752 +: 8] = op_i_flat[752 +: 8];
        op_o_flat[760 +: 8] = op_i_flat[760 +: 8];
        op_o_flat[768 +: 8] = op_i_flat[768 +: 8];
        op_o_flat[776 +: 8] = op_i_flat[776 +: 8];
        op_o_flat[784 +: 8] = op_i_flat[784 +: 8];
        op_o_flat[792 +: 8] = op_i_flat[792 +: 8];
        op_o_flat[800 +: 8] = op_i_flat[800 +: 8];
        op_o_flat[808 +: 8] = op_i_flat[808 +: 8];
        op_o_flat[816 +: 8] = op_i_flat[816 +: 8];
        op_o_flat[824 +: 8] = op_i_flat[824 +: 8];
        op_o_flat[832 +: 8] = op_i_flat[832 +: 8];
        op_o_flat[840 +: 8] = op_i_flat[840 +: 8];
        op_o_flat[848 +: 8] = op_i_flat[848 +: 8];
        op_o_flat[856 +: 8] = op_i_flat[856 +: 8];
        op_o_flat[864 +: 8] = op_i_flat[864 +: 8];
        op_o_flat[872 +: 8] = op_i_flat[872 +: 8];
        op_o_flat[880 +: 8] = op_i_flat[880 +: 8];
        op_o_flat[888 +: 8] = op_i_flat[888 +: 8];
        op_o_flat[896 +: 8] = op_i_flat[896 +: 8];
        op_o_flat[904 +: 8] = op_i_flat[904 +: 8];
        op_o_flat[912 +: 8] = op_i_flat[912 +: 8];
        op_o_flat[920 +: 8] = op_i_flat[920 +: 8];
        op_o_flat[928 +: 8] = op_i_flat[928 +: 8];
        op_o_flat[936 +: 8] = op_i_flat[936 +: 8];
        op_o_flat[944 +: 8] = op_i_flat[944 +: 8];
        op_o_flat[952 +: 8] = op_i_flat[952 +: 8];
        op_o_flat[960 +: 8] = op_i_flat[960 +: 8];
        op_o_flat[968 +: 8] = op_i_flat[968 +: 8];
        op_o_flat[976 +: 8] = op_i_flat[976 +: 8];
        op_o_flat[984 +: 8] = op_i_flat[984 +: 8];
        op_o_flat[992 +: 8] = op_i_flat[992 +: 8];
        op_o_flat[1000 +: 8] = op_i_flat[1000 +: 8];
        op_o_flat[1008 +: 8] = op_i_flat[1008 +: 8];
        op_o_flat[1016 +: 8] = op_i_flat[1016 +: 8];
      end
      default: op_o_flat = op_i_flat;
    endcase
  end
else
  $error("Error. Allowed NrLanes values are 1, 2, 4, 8, or 16");

endmodule
